CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
150 60 30 110 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
40
13 Logic Switch~
5 235 391 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6263 0 0
2
43283.1 8
0
13 Logic Switch~
5 236 453 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4900 0 0
2
43283.1 7
0
13 Logic Switch~
5 236 578 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8783 0 0
2
43283.1 6
0
13 Logic Switch~
5 235 516 0 1 11
0 23
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3221 0 0
2
43283.1 5
0
13 Logic Switch~
5 232 264 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3215 0 0
2
43283.1 1
0
13 Logic Switch~
5 233 326 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7903 0 0
2
43283.1 0
0
13 Logic Switch~
5 233 201 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7121 0 0
2
43283.1 0
0
13 Logic Switch~
5 232 139 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4484 0 0
2
43283.1 0
0
14 Logic Display~
6 811 280 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5996 0 0
2
43283.1 0
0
14 Logic Display~
6 761 280 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7804 0 0
2
43283.1 0
0
14 Logic Display~
6 717 280 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5523 0 0
2
43283.1 0
0
8 4-In OR~
219 613 380 0 5 22
0 14 7 6 5 3
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U10B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 10 0
1 U
3330 0 0
2
43283.1 0
0
8 4-In OR~
219 611 182 0 5 22
0 18 21 20 19 4
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U10A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
3465 0 0
2
43283.1 0
0
9 4-In AND~
219 501 548 0 5 22
0 10 9 8 30 2
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U9A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 9 0
1 U
8396 0 0
2
43283.1 0
0
9 2-In AND~
219 499 338 0 3 22
0 13 10 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3685 0 0
2
43283.1 2
0
5 7415~
219 500 391 0 4 22
0 12 10 9 6
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 7 0
1 U
7849 0 0
2
43283.1 1
0
9 4-In AND~
219 501 440 0 5 22
0 11 10 9 8 5
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U8B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 8 0
1 U
6343 0 0
2
43283.1 0
0
9 4-In AND~
219 499 240 0 5 22
0 15 10 9 8 19
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U8A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 8 0
1 U
7376 0 0
2
43283.1 0
0
5 7415~
219 498 191 0 4 22
0 16 10 9 20
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 7 0
1 U
9156 0 0
2
43283.1 0
0
9 2-In AND~
219 497 138 0 3 22
0 17 10 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
5776 0 0
2
43283.1 0
0
9 2-In AND~
219 328 400 0 3 22
0 34 24 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
7207 0 0
2
43283.1 13
0
9 2-In AND~
219 327 444 0 3 22
0 25 33 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
4459 0 0
2
43283.1 12
0
9 2-In NOR~
219 367 422 0 3 22
0 16 12 8
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U2D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3760 0 0
2
43283.1 11
0
5 4049~
219 283 391 0 2 22
0 25 34
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 5 0
1 U
754 0 0
2
43283.1 10
0
5 4049~
219 282 453 0 2 22
0 24 33
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 5 0
1 U
9767 0 0
2
43283.1 9
0
5 4049~
219 282 578 0 2 22
0 22 31
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 3 0
1 U
7978 0 0
2
43283.1 4
0
5 4049~
219 283 516 0 2 22
0 23 32
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 3 0
1 U
3142 0 0
2
43283.1 3
0
9 2-In NOR~
219 367 547 0 3 22
0 15 11 30
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U2C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3284 0 0
2
43283.1 2
0
9 2-In AND~
219 327 569 0 3 22
0 23 31 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
659 0 0
2
43283.1 1
0
9 2-In AND~
219 328 525 0 3 22
0 32 22 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3800 0 0
2
43283.1 0
0
9 2-In AND~
219 325 273 0 3 22
0 36 26 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
6792 0 0
2
43283.1 6
0
9 2-In AND~
219 324 317 0 3 22
0 27 35 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3701 0 0
2
43283.1 5
0
9 2-In NOR~
219 364 295 0 3 22
0 17 13 9
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
6316 0 0
2
43283.1 4
0
5 4049~
219 280 264 0 2 22
0 27 36
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
8734 0 0
2
43283.1 3
0
5 4049~
219 279 326 0 2 22
0 26 35
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
7988 0 0
2
43283.1 2
0
5 4049~
219 279 201 0 2 22
0 28 37
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
3217 0 0
2
43283.1 0
0
5 4049~
219 280 139 0 2 22
0 29 38
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
3965 0 0
2
43283.1 0
0
9 2-In NOR~
219 364 170 0 3 22
0 18 14 10
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
8239 0 0
2
43283.1 0
0
9 2-In AND~
219 324 192 0 3 22
0 29 37 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
828 0 0
2
43283.1 0
0
9 2-In AND~
219 325 148 0 3 22
0 38 28 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6187 0 0
2
43283.1 0
0
65
5 1 2 0 0 8320 0 14 11 0 0 3
522 548
717 548
717 298
5 1 3 0 0 4224 0 12 10 0 0 3
646 380
761 380
761 298
5 1 4 0 0 4224 0 13 9 0 0 5
644 182
791 182
791 306
811 306
811 298
5 4 5 0 0 4224 0 17 12 0 0 4
522 440
588 440
588 394
596 394
4 3 6 0 0 4224 0 16 12 0 0 4
521 391
588 391
588 385
596 385
3 2 7 0 0 4224 0 15 12 0 0 4
520 338
588 338
588 376
596 376
4 3 8 0 0 4096 0 17 23 0 0 4
477 454
429 454
429 422
406 422
3 3 9 0 0 8192 0 17 33 0 0 4
477 445
436 445
436 295
403 295
3 3 9 0 0 0 0 16 33 0 0 4
476 400
431 400
431 295
403 295
2 0 10 0 0 4096 0 17 0 0 41 2
477 436
411 436
2 0 10 0 0 0 0 16 0 0 41 2
476 391
411 391
2 0 10 0 0 0 0 15 0 0 41 2
475 347
411 347
3 1 11 0 0 8320 0 29 17 0 0 4
348 569
464 569
464 427
477 427
3 1 12 0 0 4224 0 22 16 0 0 4
348 444
468 444
468 382
476 382
3 1 13 0 0 4224 0 32 15 0 0 4
345 317
467 317
467 329
475 329
3 1 14 0 0 8320 0 39 12 0 0 4
345 192
470 192
470 367
596 367
4 0 8 0 0 8320 0 18 0 0 39 4
475 254
424 254
424 422
419 422
0 3 9 0 0 0 0 0 19 19 0 3
421 245
421 200
474 200
3 0 9 0 0 0 0 18 0 0 38 4
475 245
421 245
421 296
416 296
0 2 10 0 0 0 0 0 20 41 0 4
411 171
460 171
460 147
473 147
2 0 10 0 0 0 0 18 0 0 41 2
475 236
411 236
2 0 10 0 0 0 0 19 0 0 41 2
474 191
411 191
3 1 15 0 0 8320 0 30 18 0 0 4
349 525
457 525
457 227
475 227
3 1 16 0 0 8320 0 21 19 0 0 4
349 400
461 400
461 182
474 182
3 1 17 0 0 8320 0 31 20 0 0 4
346 273
465 273
465 129
473 129
3 1 18 0 0 12416 0 40 13 0 0 4
346 148
469 148
469 169
594 169
5 4 19 0 0 4224 0 18 13 0 0 4
520 240
586 240
586 196
594 196
4 3 20 0 0 4224 0 19 13 0 0 4
519 191
586 191
586 187
594 187
3 2 21 0 0 4224 0 20 13 0 0 4
518 138
586 138
586 178
594 178
1 2 22 0 0 12416 0 26 30 0 0 4
267 578
258 578
258 534
304 534
1 1 23 0 0 8320 0 27 29 0 0 4
268 516
264 516
264 560
303 560
1 2 24 0 0 12416 0 25 21 0 0 4
267 453
258 453
258 409
304 409
1 1 25 0 0 8320 0 24 22 0 0 4
268 391
264 391
264 435
303 435
1 2 26 0 0 12416 0 35 31 0 0 4
264 326
255 326
255 282
301 282
1 1 27 0 0 8320 0 34 32 0 0 4
265 264
261 264
261 308
300 308
1 2 28 0 0 12416 0 36 40 0 0 4
264 201
255 201
255 157
301 157
1 1 29 0 0 8320 0 37 39 0 0 4
265 139
261 139
261 183
300 183
2 3 9 0 0 8320 0 14 33 0 0 4
477 544
416 544
416 295
403 295
3 3 8 0 0 128 0 14 23 0 0 4
477 553
419 553
419 422
406 422
4 3 30 0 0 4224 0 14 28 0 0 4
477 562
414 562
414 547
406 547
1 3 10 0 0 8320 0 14 38 0 0 4
477 535
411 535
411 170
403 170
1 1 22 0 0 0 0 3 26 0 0 2
248 578
267 578
1 1 23 0 0 0 0 4 27 0 0 2
247 516
268 516
2 2 31 0 0 0 0 26 29 0 0 2
303 578
303 578
2 1 32 0 0 0 0 27 30 0 0 2
304 516
304 516
3 2 11 0 0 128 0 29 28 0 0 3
348 569
348 556
354 556
3 1 15 0 0 128 0 30 28 0 0 3
349 525
349 538
354 538
1 1 24 0 0 0 0 2 25 0 0 2
248 453
267 453
1 1 25 0 0 0 0 1 24 0 0 2
247 391
268 391
2 2 33 0 0 0 0 25 22 0 0 2
303 453
303 453
2 1 34 0 0 0 0 24 21 0 0 2
304 391
304 391
3 2 12 0 0 128 0 22 23 0 0 3
348 444
348 431
354 431
3 1 16 0 0 128 0 21 23 0 0 3
349 400
349 413
354 413
1 1 26 0 0 0 0 6 35 0 0 2
245 326
264 326
1 1 27 0 0 0 0 5 34 0 0 2
244 264
265 264
2 2 35 0 0 0 0 35 32 0 0 2
300 326
300 326
2 1 36 0 0 0 0 34 31 0 0 2
301 264
301 264
3 2 13 0 0 128 0 32 33 0 0 3
345 317
345 304
351 304
3 1 17 0 0 128 0 31 33 0 0 3
346 273
346 286
351 286
1 1 28 0 0 0 0 7 36 0 0 2
245 201
264 201
1 1 29 0 0 0 0 8 37 0 0 2
244 139
265 139
2 2 37 0 0 0 0 36 39 0 0 2
300 201
300 201
2 1 38 0 0 0 0 37 40 0 0 2
301 139
301 139
3 2 14 0 0 128 0 39 38 0 0 3
345 192
345 179
351 179
3 1 18 0 0 128 0 40 38 0 0 3
346 148
346 161
351 161
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
788 233 831 255
797 241 821 257
3 A<B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
738 234 781 256
747 241 771 257
3 A>B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
695 234 738 256
704 241 728 257
3 A=B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
381 144 414 165
389 151 405 166
2 X3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
379 268 414 289
388 275 404 290
2 X2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
383 394 418 415
392 401 408 416
2 X1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
385 519 418 540
393 525 409 540
2 X0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
