CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
208 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
376 176 489 273
9437202 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 304 333 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 ONE
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43283.1 0
0
13 Logic Switch~
5 299 245 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
43283.1 1
0
13 Logic Switch~
5 300 279 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
43283.1 0
0
13 Logic Switch~
5 300 210 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
43283.1 0
0
13 Logic Switch~
5 302 145 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
43283.1 0
0
14 Logic Display~
6 554 245 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
43283.1 0
0
9 Inverter~
13 350 145 0 2 22
0 4 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
8901 0 0
2
43283.1 0
0
9 Inverter~
13 355 333 0 2 22
0 6 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
7361 0 0
2
43283.1 0
0
6 CD4512
77 442 241 0 14 29
0 4 3 3 5 5 3 6 6 9
8 7 3 3 2
0
0 0 4336 0
4 4512
-14 -60 14 -52
2 U1
-7 -70 7 -62
0
15 DVDD=16;DGND=8;
146 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 7 6 5 4 3 2 1 13
12 11 15 10 14 9 7 6 5 4
3 2 1 13 12 11 15 10 14 0
65 0 0 0 0 0 0 0
1 U
4747 0 0
2
43283.1 0
0
16
14 1 2 0 0 4240 0 9 6 0 0 3
474 277
554 277
554 263
12 0 3 0 0 4096 0 9 0 0 3 2
480 250
499 250
13 0 3 0 0 12416 0 9 0 0 12 6
480 259
499 259
499 170
387 170
387 223
397 223
0 1 4 0 0 8320 0 0 9 7 0 3
330 145
330 214
410 214
4 0 5 0 0 4096 0 9 0 0 6 2
410 241
392 241
2 5 5 0 0 8320 0 7 9 0 0 4
371 145
392 145
392 250
410 250
1 1 4 0 0 0 0 5 7 0 0 2
314 145
335 145
0 8 6 0 0 4096 0 0 9 9 0 3
405 268
405 277
410 277
0 7 6 0 0 8320 0 0 9 13 0 3
327 333
327 268
410 268
0 6 3 0 0 0 0 0 9 12 0 2
397 259
410 259
0 3 3 0 0 0 0 0 9 12 0 2
397 232
410 232
2 2 3 0 0 128 0 8 9 0 0 4
376 333
397 333
397 223
410 223
1 1 6 0 0 0 0 1 8 0 0 2
316 333
340 333
1 11 7 0 0 8320 0 3 9 0 0 6
312 279
401 279
401 175
493 175
493 232
474 232
1 10 8 0 0 4224 0 2 9 0 0 6
311 245
406 245
406 180
488 180
488 223
474 223
9 1 9 0 0 12416 0 9 4 0 0 6
474 214
484 214
484 185
323 185
323 210
312 210
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
