CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 501 178 0 1 11
0 9
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4722 0 0
2
5.89748e-315 0
0
13 Logic Switch~
5 122 348 0 1 11
0 16
0
0 0 21344 0
2 0V
-30 0 -16 8
2 V9
-29 -10 -15 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
386 0 0
2
5.89748e-315 0
0
13 Logic Switch~
5 122 316 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-31 -1 -17 7
2 V8
-31 -14 -17 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3141 0 0
2
5.89748e-315 0
0
13 Logic Switch~
5 124 285 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-31 0 -17 8
2 V7
-32 -13 -18 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3191 0 0
2
5.89748e-315 0
0
13 Logic Switch~
5 124 256 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-30 -1 -16 7
2 V6
-30 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3488 0 0
2
5.89748e-315 0
0
13 Logic Switch~
5 124 226 0 1 11
0 20
0
0 0 21344 0
2 0V
-31 -2 -17 6
2 V5
-32 -12 -18 -4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7538 0 0
2
5.89748e-315 0
0
13 Logic Switch~
5 125 201 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-31 0 -17 8
2 V4
-30 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3386 0 0
2
5.89748e-315 0
0
13 Logic Switch~
5 125 175 0 1 11
0 22
0
0 0 21344 0
2 0V
-33 0 -19 8
2 V3
-32 -11 -18 -3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3249 0 0
2
5.89748e-315 0
0
13 Logic Switch~
5 125 149 0 1 11
0 23
0
0 0 21344 0
2 0V
-28 0 -14 8
2 V2
-28 -13 -14 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
374 0 0
2
5.89748e-315 0
0
13 Logic Switch~
5 123 125 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-31 0 -17 8
2 V1
-31 -12 -17 -4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3579 0 0
2
5.89748e-315 0
0
14 Logic Display~
6 437 177 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
871 0 0
2
5.89748e-315 0
0
14 Logic Display~
6 796 133 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
985 0 0
2
5.89748e-315 0
0
14 Logic Display~
6 775 135 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5843 0 0
2
5.89748e-315 0
0
14 Logic Display~
6 755 135 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7221 0 0
2
5.89748e-315 0
0
14 Logic Display~
6 732 138 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6830 0 0
2
5.89748e-315 0
0
14 Logic Display~
6 709 139 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3945 0 0
2
5.89748e-315 0
0
8 3-In OR~
219 503 113 0 4 22
0 11 10 3 2
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 3 0
1 U
4623 0 0
2
5.89748e-315 0
0
9 2-In AND~
219 405 76 0 3 22
0 13 14 11
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
8115 0 0
2
5.89748e-315 0
0
5 4081~
219 414 149 0 3 22
0 13 12 10
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
360 0 0
2
5.89748e-315 0
0
4 4008
219 651 215 0 14 29
0 9 2 2 9 13 14 12 15 2
4 5 6 7 8
0
0 0 4832 0
4 4008
-14 -60 14 -52
2 U2
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 0 1 0 0 0
1 U
3628 0 0
2
5.89748e-315 0
0
4 4008
219 312 232 0 14 29
0 24 23 22 21 20 19 18 17 16
15 12 14 13 3
0
0 0 4832 0
4 4008
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 0 1 0 0 0
1 U
7221 0 0
2
5.89748e-315 0
0
31
0 9 2 0 0 4224 0 0 20 11 0 3
556 113
556 251
619 251
1 0 3 0 0 4096 0 11 0 0 12 2
437 195
437 196
10 1 4 0 0 4224 0 20 12 0 0 3
683 224
796 224
796 151
11 1 5 0 0 4224 0 20 13 0 0 3
683 215
775 215
775 153
12 1 6 0 0 4224 0 20 14 0 0 3
683 206
755 206
755 153
13 1 7 0 0 4224 0 20 15 0 0 3
683 197
732 197
732 156
14 1 8 0 0 4224 0 20 16 0 0 3
683 179
709 179
709 157
0 4 9 0 0 8192 0 0 20 9 0 3
548 178
548 206
619 206
1 1 9 0 0 4224 0 1 20 0 0 4
513 178
606 178
606 179
619 179
0 3 2 0 0 0 0 0 20 11 0 3
611 188
611 197
619 197
4 2 2 0 0 0 0 17 20 0 0 4
536 113
611 113
611 188
619 188
14 3 3 0 0 4224 0 21 17 0 0 4
344 196
477 196
477 122
490 122
3 2 10 0 0 4224 0 19 17 0 0 4
435 149
484 149
484 113
491 113
3 1 11 0 0 4224 0 18 17 0 0 4
426 76
484 76
484 104
490 104
0 2 12 0 0 4096 0 0 19 21 0 3
380 232
380 158
390 158
0 1 13 0 0 4096 0 0 19 18 0 2
370 140
390 140
0 2 14 0 0 4096 0 0 18 20 0 3
361 223
361 85
381 85
0 1 13 0 0 4096 0 0 18 19 0 3
370 214
370 67
381 67
13 5 13 0 0 12416 0 21 20 0 0 4
344 214
370 214
370 215
619 215
12 6 14 0 0 12416 0 21 20 0 0 4
344 223
361 223
361 224
619 224
11 7 12 0 0 12416 0 21 20 0 0 4
344 232
380 232
380 233
619 233
10 8 15 0 0 12416 0 21 20 0 0 4
344 241
359 241
359 242
619 242
1 9 16 0 0 4224 0 2 21 0 0 4
134 348
262 348
262 268
280 268
1 8 17 0 0 4224 0 3 21 0 0 4
134 316
272 316
272 259
280 259
1 7 18 0 0 4224 0 4 21 0 0 4
136 285
266 285
266 250
280 250
1 6 19 0 0 4224 0 5 21 0 0 4
136 256
254 256
254 241
280 241
1 5 20 0 0 4224 0 6 21 0 0 4
136 226
259 226
259 232
280 232
1 4 21 0 0 4224 0 7 21 0 0 4
137 201
259 201
259 223
280 223
1 3 22 0 0 4224 0 8 21 0 0 4
137 175
249 175
249 214
280 214
1 2 23 0 0 4224 0 9 21 0 0 4
137 149
254 149
254 205
280 205
1 1 24 0 0 4224 0 10 21 0 0 4
135 125
259 125
259 196
280 196
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
