CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
6
13 Logic Switch~
5 200 201 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-10 12 4 20
1 B
-25 -1 -18 7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
42398.9 0
0
13 Logic Switch~
5 203 179 0 1 11
0 5
0
0 0 21344 0
2 0V
-10 -20 4 -12
1 A
-27 -4 -20 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.8974e-315 0
0
14 Logic Display~
6 597 253 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3124 0 0
2
5.8974e-315 0
0
14 Logic Display~
6 604 175 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3421 0 0
2
5.8974e-315 0
0
5 4081~
219 440 271 0 3 22
0 5 4 2
0
0 0 96 0
4 4081
-7 -24 21 -16
2 A1
0 -34 14 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
8157 0 0
2
5.8974e-315 0
0
5 4030~
219 429 188 0 3 22
0 5 4 3
0
0 0 96 0
4 4030
-7 -24 21 -16
2 A2
0 -34 14 -26
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
5572 0 0
2
5.8974e-315 0
0
6
1 2 0 0 0 0 0 1 6 0 0 4
212 201
405 201
405 197
413 197
3 1 2 0 0 4224 0 5 3 0 0 2
461 271
597 271
3 1 3 0 0 4224 0 6 4 0 0 3
462 188
604 188
604 193
0 2 4 0 0 4096 0 0 5 0 0 3
354 205
354 280
416 280
0 1 5 0 0 8192 0 0 5 6 0 3
319 179
319 262
416 262
1 1 5 0 0 4224 0 2 6 0 0 2
215 179
413 179
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
343 331 442 352
352 338 432 353
10 Half Adder
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
508 173 551 194
517 179 541 194
3 SUM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
478 250 537 271
487 257 527 272
5 CARRY
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
