CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 151 39 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 G3
-30 0 -16 8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3820 0 0
2
42398.9 18
0
13 Logic Switch~
5 153 170 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 P3
-29 -1 -15 7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7678 0 0
2
42398.9 17
0
13 Logic Switch~
5 162 354 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 P2
-30 -2 -16 6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
961 0 0
2
42398.9 16
0
13 Logic Switch~
5 159 270 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 G2
-30 -5 -16 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3178 0 0
2
42398.9 15
0
13 Logic Switch~
5 162 423 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 G1
-29 -3 -15 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3409 0 0
2
42398.9 14
0
13 Logic Switch~
5 165 461 0 1 11
0 13
0
0 0 21360 0
2 0V
-5 -17 9 -9
2 P1
-32 0 -18 8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3951 0 0
2
42398.9 13
0
13 Logic Switch~
5 165 509 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 C1
-34 -2 -20 6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8885 0 0
2
42398.9 12
0
14 Logic Display~
6 1054 474 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3780 0 0
2
42398.9 11
0
14 Logic Display~
6 1058 291 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9265 0 0
2
42398.9 10
0
14 Logic Display~
6 1053 113 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9442 0 0
2
42398.9 9
0
8 4-In OR~
219 787 132 0 5 22
0 8 7 6 5 4
0
0 0 112 0
4 4072
-14 -24 14 -16
0
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
9424 0 0
2
42398.9 8
0
5 4081~
219 516 94 0 3 22
0 10 9 7
0
0 0 112 0
4 4081
-7 -24 21 -16
0
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
9968 0 0
2
42398.9 7
0
5 4073~
219 517 137 0 4 22
0 10 12 11 6
0
0 0 112 0
4 4073
-7 -24 21 -16
0
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 3 0
1 U
9281 0 0
2
42398.9 6
0
5 4082~
219 517 186 0 5 22
0 10 12 13 14 5
0
0 0 112 0
4 4082
-7 -24 21 -16
0
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
8464 0 0
2
42398.9 5
0
8 3-In OR~
219 785 308 0 4 22
0 9 15 16 3
0
0 0 112 0
4 4075
-14 -24 14 -16
0
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
7168 0 0
2
42398.9 4
0
5 4081~
219 516 308 0 3 22
0 12 11 15
0
0 0 112 0
4 4081
-7 -24 21 -16
0
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
3171 0 0
2
42398.9 3
0
5 4073~
219 517 364 0 4 22
0 12 13 14 16
0
0 0 112 0
4 4073
-7 -24 21 -16
0
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 3 0
1 U
4139 0 0
2
42398.9 2
0
5 4071~
219 791 491 0 3 22
0 11 17 2
0
0 0 112 0
4 4071
-7 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
6435 0 0
2
42398.9 1
0
5 4081~
219 519 500 0 3 22
0 13 14 17
0
0 0 112 0
4 4081
-7 -24 21 -16
0
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
5283 0 0
2
42398.9 0
0
28
3 1 2 0 0 4240 0 18 8 0 0 3
824 491
1054 491
1054 492
4 1 3 0 0 4240 0 15 9 0 0 3
818 308
1058 308
1058 309
5 1 4 0 0 4240 0 11 10 0 0 3
820 132
1053 132
1053 131
5 4 5 0 0 12432 0 14 11 0 0 4
538 186
553 186
553 146
770 146
4 3 6 0 0 4240 0 13 11 0 0 2
538 137
770 137
3 2 7 0 0 4240 0 12 11 0 0 4
537 94
754 94
754 128
770 128
1 1 8 0 0 4240 0 1 11 0 0 4
163 39
759 39
759 119
770 119
0 2 9 0 0 4112 0 0 12 17 0 3
330 270
330 103
492 103
0 1 10 0 0 8208 0 0 12 12 0 3
246 128
246 85
492 85
0 3 11 0 0 4112 0 0 13 21 0 3
407 317
407 146
493 146
0 2 12 0 0 8208 0 0 13 13 0 3
289 182
289 137
493 137
0 1 10 0 0 8208 0 0 13 16 0 3
212 170
212 128
493 128
0 2 12 0 0 8208 0 0 14 20 0 3
257 299
257 182
493 182
0 3 13 0 0 4112 0 0 14 22 0 3
376 364
376 191
493 191
0 4 14 0 0 4112 0 0 14 24 0 3
460 373
460 200
493 200
1 1 10 0 0 4240 0 2 14 0 0 4
165 170
485 170
485 173
493 173
1 1 9 0 0 4240 0 4 15 0 0 4
171 270
763 270
763 299
772 299
3 2 15 0 0 4240 0 16 15 0 0 2
537 308
773 308
4 3 16 0 0 4240 0 17 15 0 0 4
538 364
763 364
763 317
772 317
0 1 12 0 0 8208 0 0 16 23 0 3
240 354
240 299
492 299
0 2 11 0 0 16 0 0 16 25 0 3
348 423
348 317
492 317
0 2 13 0 0 8208 0 0 17 28 0 3
211 461
211 364
493 364
1 1 12 0 0 4240 0 3 17 0 0 4
174 354
472 354
472 355
493 355
0 3 14 0 0 16 0 0 17 27 0 3
393 509
393 373
493 373
1 1 11 0 0 4240 0 5 18 0 0 4
174 423
768 423
768 482
778 482
3 2 17 0 0 4240 0 19 18 0 0 2
540 500
778 500
1 2 14 0 0 4240 0 7 19 0 0 2
177 509
495 509
1 1 13 0 0 4240 0 6 19 0 0 4
177 461
492 461
492 491
495 491
11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
467 552 560 576
477 560 549 576
9 Generator
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
329 550 478 574
339 558 467 574
16 Look Ahead Carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
867 460 904 484
877 468 893 484
2 C2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
857 284 902 308
867 292 891 308
3  C3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
830 108 907 132
840 116 896 132
7      C4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
608 69 661 93
618 77 650 93
4 P3G2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
610 110 679 134
620 118 668 134
6 P3P2G1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
610 145 695 169
620 153 684 169
8 P3P2P1C1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
582 283 635 307
592 291 624 307
4 G1P2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
579 338 648 362
589 346 637 362
6 P2P1C1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
598 475 651 499
608 483 640 499
4 P1C1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
