CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 110 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 89 350 0 1 11
0 6
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 Cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.8974e-315 0
0
13 Logic Switch~
5 83 177 0 1 11
0 8
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.8974e-315 0
0
13 Logic Switch~
5 148 147 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.8974e-315 0
0
14 Logic Display~
6 1019 262 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3421 0 0
2
5.8974e-315 0
0
14 Logic Display~
6 863 157 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.8974e-315 0
0
5 4071~
219 880 279 0 3 22
0 4 5 2
0
0 0 96 0
4 4071
-7 -24 21 -16
2 A1
0 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
5572 0 0
2
5.8974e-315 0
0
5 4081~
219 669 290 0 3 22
0 7 6 5
0
0 0 96 0
4 4081
-7 -24 21 -16
2 A2
0 -34 14 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
8901 0 0
2
5.8974e-315 0
0
5 4081~
219 417 235 0 3 22
0 9 8 4
0
0 0 96 0
4 4081
-7 -24 21 -16
2 A3
0 -34 14 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
7361 0 0
2
5.8974e-315 0
0
5 4070~
219 653 174 0 3 22
0 7 6 3
0
0 0 96 0
4 4070
-7 -24 21 -16
2 A4
0 -34 14 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
4747 0 0
2
5.8974e-315 0
0
5 4070~
219 400 164 0 3 22
0 9 8 7
0
0 0 96 0
4 4070
-7 -24 21 -16
2 A5
0 -34 14 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
972 0 0
2
5.8974e-315 0
0
12
3 1 2 0 0 4224 0 6 4 0 0 3
913 279
1019 279
1019 280
3 1 3 0 0 4224 0 9 5 0 0 3
686 174
863 174
863 175
3 1 4 0 0 4224 0 8 6 0 0 4
438 235
859 235
859 270
867 270
3 2 5 0 0 4224 0 7 6 0 0 4
690 290
859 290
859 288
867 288
0 2 6 0 0 4096 0 0 7 7 0 2
607 299
645 299
0 1 7 0 0 4096 0 0 7 8 0 3
561 165
561 281
645 281
1 2 6 0 0 4224 0 1 9 0 0 4
101 350
607 350
607 183
637 183
3 1 7 0 0 12416 0 10 9 0 0 4
433 164
448 164
448 165
637 165
0 2 8 0 0 8192 0 0 8 11 0 3
310 177
310 244
393 244
0 1 9 0 0 8192 0 0 8 12 0 3
262 147
262 226
393 226
1 2 8 0 0 4224 0 2 10 0 0 4
95 177
376 177
376 173
384 173
1 1 9 0 0 4224 0 3 10 0 0 4
160 147
376 147
376 155
384 155
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
299 392 398 414
308 399 388 415
10 Full Adder
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
713 147 758 171
723 155 747 171
3 SUM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
938 255 999 279
948 263 988 279
5 CARRY
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
