CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
390 170 30 400 10
176 79 1358 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 426 232 0 1 11
0 11
0
0 0 21360 0
2 0V
-29 -2 -15 6
2 V4
-27 -11 -13 -3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
42461 0
0
13 Logic Switch~
5 425 297 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-29 1 -15 9
2 V3
-28 -8 -14 0
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
42461 0
0
13 Logic Switch~
5 425 274 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-29 -3 -15 5
2 V2
-29 -12 -15 -4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
42461 0
0
13 Logic Switch~
5 425 253 0 1 11
0 12
0
0 0 21360 0
2 0V
-29 -1 -15 7
2 V1
-29 -12 -15 -4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
42461 0
0
14 Logic Display~
6 669 272 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
42461 0
0
14 Logic Display~
6 667 213 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
42461 0
0
8 4-In OR~
219 621 290 0 5 22
0 4 8 9 10 2
0
0 0 624 0
4 4072
-14 -24 14 -16
1 S
4 -25 11 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 1 0
1 U
8901 0 0
2
42461 0
0
8 4-In OR~
219 615 232 0 5 22
0 4 5 6 7 3
0
0 0 624 0
4 4072
-14 -24 14 -16
4 Cout
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 1 0
1 U
7361 0 0
2
42461 0
0
4 4028
219 522 253 0 14 29
0 11 12 13 14 15 10 9 7 8
6 5 4 16 17
0
0 0 4848 0
4 4028
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
106 %D [%16bi %8bi %1i %2i %3i %4i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 12 13 10 3 14 2 15 1
6 7 4 9 5 11 12 13 10 3
14 2 15 1 6 7 4 9 5 0
65 0 0 512 0 0 0 0
1 U
4747 0 0
2
42461 0
0
14
5 1 2 0 0 4224 0 7 5 0 0 2
654 290
669 290
5 1 3 0 0 12416 0 8 6 0 0 5
648 232
655 232
655 239
667 239
667 231
0 1 4 0 0 8192 0 0 8 7 0 3
569 235
569 219
598 219
11 2 5 0 0 4224 0 9 8 0 0 4
554 244
585 244
585 228
598 228
10 3 6 0 0 4224 0 9 8 0 0 4
554 253
580 253
580 237
598 237
8 4 7 0 0 4224 0 9 8 0 0 4
554 271
585 271
585 246
598 246
12 1 4 0 0 8320 0 9 7 0 0 4
554 235
589 235
589 277
604 277
9 2 8 0 0 4224 0 9 7 0 0 4
554 262
596 262
596 286
604 286
7 3 9 0 0 4224 0 9 7 0 0 4
554 280
591 280
591 295
604 295
6 4 10 0 0 4224 0 9 7 0 0 4
554 289
596 289
596 304
604 304
1 1 11 0 0 4224 0 1 9 0 0 4
438 232
482 232
482 271
490 271
1 2 12 0 0 4224 0 4 9 0 0 4
437 253
477 253
477 280
490 280
1 3 13 0 0 4224 0 3 9 0 0 4
437 274
482 274
482 289
490 289
1 4 14 0 0 4224 0 2 9 0 0 4
437 297
482 297
482 298
490 298
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
