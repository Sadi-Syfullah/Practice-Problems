CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
80 10 30 150 10
176 79 1358 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
16
13 Logic Switch~
5 241 262 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
42469 0
0
13 Logic Switch~
5 241 227 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
42469 0
0
13 Logic Switch~
5 241 191 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
42469 0
0
13 Logic Switch~
5 242 152 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
42469 0
0
5 7422~
219 727 275 0 5 22
0 10 12 13 11 2
0
0 0 624 0
6 74LS22
-21 -28 21 -20
3 U4B
-12 -31 9 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 3 0
1 U
8157 0 0
2
42469 0
0
5 7422~
219 731 115 0 5 22
0 6 4 5 10 3
0
0 0 624 0
6 74LS22
-21 -28 21 -20
3 U4A
-12 -31 9 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 3 0
1 U
5572 0 0
2
42469 0
0
10 2-In NAND~
219 591 367 0 3 22
0 17 17 11
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
8901 0 0
2
42469 0
0
10 2-In NAND~
219 588 43 0 3 22
0 7 7 6
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7361 0 0
2
42469 0
0
10 2-In NAND~
219 589 317 0 3 22
0 16 16 12
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
4747 0 0
2
42469 0
0
10 2-In NAND~
219 585 259 0 3 22
0 15 15 13
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
972 0 0
2
42469 0
0
10 2-In NAND~
219 585 197 0 3 22
0 14 14 10
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3472 0 0
2
42469 0
0
10 2-In NAND~
219 584 149 0 3 22
0 9 9 4
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9998 0 0
2
42469 0
0
10 2-In NAND~
219 586 94 0 3 22
0 8 8 5
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3536 0 0
2
42469 0
0
14 Logic Display~
6 828 219 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4597 0 0
2
42469 0
0
14 Logic Display~
6 823 119 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3835 0 0
2
42469 0
0
4 4028
219 421 189 0 14 29
0 18 19 20 21 22 17 16 9 15
8 7 14 23 24
0
0 0 4848 0
4 4028
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
106 %D [%16bi %8bi %1i %2i %3i %4i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 12 13 10 3 14 2 15 1
6 7 4 9 5 11 12 13 10 3
14 2 15 1 6 7 4 9 5 0
65 0 0 512 0 0 0 0
1 U
3670 0 0
2
42469 0
0
28
5 1 2 0 0 4224 0 5 14 0 0 3
754 275
828 275
828 237
5 1 3 0 0 4224 0 6 15 0 0 5
758 115
811 115
811 145
823 145
823 137
3 2 4 0 0 4224 0 12 6 0 0 4
611 149
699 149
699 121
707 121
3 3 5 0 0 4224 0 13 6 0 0 4
613 94
694 94
694 109
707 109
3 1 6 0 0 4224 0 8 6 0 0 4
615 43
699 43
699 97
707 97
0 2 7 0 0 8192 0 0 8 7 0 3
556 53
556 52
564 52
11 1 7 0 0 8320 0 16 8 0 0 4
453 180
556 180
556 34
564 34
0 1 8 0 0 4096 0 0 13 9 0 3
552 103
552 85
562 85
10 2 8 0 0 4224 0 16 13 0 0 4
453 189
539 189
539 103
562 103
0 2 9 0 0 4096 0 0 12 11 0 3
547 140
547 158
560 158
8 1 9 0 0 4224 0 16 12 0 0 4
453 207
542 207
542 140
560 140
0 4 10 0 0 8192 0 0 6 16 0 3
629 197
629 133
707 133
3 4 11 0 0 8320 0 7 5 0 0 4
618 367
690 367
690 293
703 293
3 2 12 0 0 4224 0 9 5 0 0 4
616 317
695 317
695 281
703 281
3 3 13 0 0 4224 0 10 5 0 0 4
612 259
695 259
695 269
703 269
3 1 10 0 0 4224 0 11 5 0 0 4
612 197
695 197
695 257
703 257
0 2 14 0 0 4096 0 0 11 18 0 3
553 187
553 206
561 206
12 1 14 0 0 4224 0 16 11 0 0 4
453 171
553 171
553 188
561 188
0 2 15 0 0 8192 0 0 10 20 0 4
548 249
543 249
543 268
561 268
9 1 15 0 0 4224 0 16 10 0 0 4
453 198
548 198
548 250
561 250
0 2 16 0 0 8192 0 0 9 22 0 4
552 308
547 308
547 326
565 326
7 1 16 0 0 4224 0 16 9 0 0 4
453 216
552 216
552 308
565 308
0 2 17 0 0 8192 0 0 7 24 0 4
556 357
559 357
559 376
567 376
6 1 17 0 0 8320 0 16 7 0 0 4
453 225
556 225
556 358
567 358
1 1 18 0 0 4224 0 4 16 0 0 4
254 152
376 152
376 207
389 207
1 2 19 0 0 4224 0 3 16 0 0 4
253 191
381 191
381 216
389 216
1 3 20 0 0 4224 0 2 16 0 0 4
253 227
381 227
381 225
389 225
1 4 21 0 0 4224 0 1 16 0 0 4
253 262
381 262
381 234
389 234
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
