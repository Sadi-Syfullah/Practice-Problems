CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 237 86 0 1 11
0 23
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 Cin
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89852e-315 0
0
13 Logic Switch~
5 475 38 0 1 11
0 11
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89852e-315 5.32571e-315
0
13 Logic Switch~
5 460 38 0 1 11
0 12
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89852e-315 5.30499e-315
0
13 Logic Switch~
5 443 37 0 1 11
0 13
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89852e-315 5.26354e-315
0
13 Logic Switch~
5 426 37 0 1 11
0 14
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.89852e-315 0
0
13 Logic Switch~
5 383 36 0 1 11
0 15
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.89852e-315 5.32571e-315
0
13 Logic Switch~
5 367 36 0 1 11
0 16
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.89852e-315 5.30499e-315
0
13 Logic Switch~
5 351 36 0 1 11
0 17
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
5.89852e-315 5.26354e-315
0
13 Logic Switch~
5 332 36 0 1 11
0 18
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
5.89852e-315 0
0
13 Logic Switch~
5 236 314 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
5.89852e-315 0
0
8 2-In OR~
219 325 413 0 3 22
0 6 2 5
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U5A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3472 0 0
2
5.89852e-315 0
0
14 Logic Display~
6 587 358 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
5.89852e-315 0
0
8 3-In OR~
219 268 266 0 4 22
0 3 21 2 22
0
0 0 624 270
4 4075
-14 -24 14 -16
3 U4A
28 -7 49 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
3536 0 0
2
5.89852e-315 0
0
9 2-In AND~
219 337 248 0 3 22
0 19 4 3
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U3B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
4597 0 0
2
5.89852e-315 0
0
9 2-In AND~
219 336 205 0 3 22
0 20 4 21
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U3A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3835 0 0
2
5.89852e-315 0
0
14 Logic Display~
6 477 357 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Carry
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
5.89852e-315 5.26354e-315
0
14 Logic Display~
6 508 358 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
5.89852e-315 0
0
14 Logic Display~
6 534 358 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
5.89852e-315 0
0
14 Logic Display~
6 561 358 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
5.89852e-315 0
0
7 74LS283
152 380 357 0 14 29
0 4 20 19 25 24 22 22 24 24
7 8 9 10 6
0
0 0 4848 270
6 74F283
-21 -60 21 -52
2 U2
57 -2 71 6
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 0 1 0 0 0
1 U
3108 0 0
2
5.89852e-315 0
0
7 74LS283
152 385 119 0 14 29
0 14 13 12 11 18 17 16 15 23
4 20 19 25 2
0
0 0 4848 270
6 74F283
-21 -60 21 -52
2 U1
57 -2 71 6
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 0 1 0 0 0
1 U
4299 0 0
2
5.89852e-315 0
0
32
0 2 2 0 0 4224 0 0 11 4 0 4
307 186
307 382
319 382
319 397
3 1 3 0 0 12416 0 14 13 0 0 5
310 248
297 248
297 235
280 235
280 250
2 0 4 0 0 4096 0 15 0 0 32 2
354 196
396 196
14 3 2 0 0 0 0 21 13 0 0 4
342 153
342 186
262 186
262 250
3 1 5 0 0 4224 0 11 16 0 0 3
328 443
477 443
477 375
14 1 6 0 0 4224 0 20 11 0 0 2
337 391
337 397
10 1 7 0 0 8320 0 20 17 0 0 4
391 391
391 410
508 410
508 376
11 1 8 0 0 8320 0 20 18 0 0 4
382 391
382 405
534 405
534 376
12 1 9 0 0 8320 0 20 19 0 0 4
373 391
373 400
561 400
561 376
13 1 10 0 0 8320 0 20 12 0 0 4
364 391
364 395
587 395
587 376
1 4 11 0 0 8320 0 2 21 0 0 4
475 50
475 66
396 66
396 89
1 3 12 0 0 8320 0 3 21 0 0 4
460 50
460 71
405 71
405 89
1 2 13 0 0 8320 0 4 21 0 0 4
443 49
443 76
414 76
414 89
1 1 14 0 0 4224 0 5 21 0 0 4
426 49
426 81
423 81
423 89
1 8 15 0 0 8320 0 6 21 0 0 4
383 48
383 66
360 66
360 89
1 7 16 0 0 4224 0 7 21 0 0 4
367 48
367 71
369 71
369 89
1 6 17 0 0 4224 0 8 21 0 0 4
351 48
351 76
378 76
378 89
1 5 18 0 0 8320 0 9 21 0 0 4
332 48
332 81
387 81
387 89
1 0 19 0 0 4096 0 14 0 0 30 2
355 257
378 257
2 0 4 0 0 0 0 14 0 0 32 2
355 239
396 239
1 0 20 0 0 4096 0 15 0 0 31 2
354 214
387 214
3 2 21 0 0 8320 0 15 13 0 0 3
309 205
271 205
271 251
7 0 22 0 0 4096 0 20 0 0 24 2
364 327
364 309
4 6 22 0 0 8320 0 13 20 0 0 4
271 296
271 309
373 309
373 327
1 9 23 0 0 4224 0 1 21 0 0 3
249 86
342 86
342 89
0 9 24 0 0 4096 0 0 20 28 0 2
337 314
337 327
8 0 24 0 0 0 0 20 0 0 28 2
355 327
355 314
1 5 24 0 0 4224 0 10 20 0 0 3
248 314
382 314
382 327
13 4 25 0 0 4224 0 21 20 0 0 4
369 153
369 319
391 319
391 327
12 3 19 0 0 4224 0 21 20 0 0 4
378 153
378 309
400 309
400 327
11 2 20 0 0 4224 0 21 20 0 0 4
387 153
387 314
409 314
409 327
10 1 4 0 0 4224 0 21 20 0 0 4
396 153
396 319
418 319
418 327
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
