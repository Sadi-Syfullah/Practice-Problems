CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
280 130 30 200 10
176 79 1358 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 362 331 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-28 -2 -14 6
2 V6
-28 -13 -14 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
42460.9 0
0
13 Logic Switch~
5 361 304 0 1 11
0 2
0
0 0 21360 0
2 0V
-30 2 -16 10
2 V5
-28 -9 -14 -1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
42460.9 0
0
13 Logic Switch~
5 361 277 0 1 11
0 9
0
0 0 21360 0
2 0V
-31 0 -17 8
2 V4
-30 -11 -16 -3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
42460.9 0
0
13 Logic Switch~
5 363 257 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-31 0 -17 8
2 V3
-30 -11 -16 -3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
42460.9 0
0
13 Logic Switch~
5 362 229 0 1 11
0 10
0
0 0 21360 0
2 0V
-34 -1 -20 7
2 V2
-33 -12 -19 -4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8157 0 0
2
42460.9 0
0
13 Logic Switch~
5 363 205 0 1 11
0 11
0
0 0 21360 0
2 0V
-34 0 -20 8
2 V1
-32 -12 -18 -4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5572 0 0
2
42460.9 0
0
14 Logic Display~
6 689 214 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
42460.9 0
0
14 Logic Display~
6 731 235 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7361 0 0
2
42460.9 0
0
14 Logic Display~
6 773 249 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
42460.9 0
0
14 Logic Display~
6 811 265 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
972 0 0
2
42460.9 0
0
4 4008
219 518 279 0 14 29
0 11 10 8 9 2 2 7 7 2
6 5 4 3 12
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 0 0 0 0
1 U
3472 0 0
2
42460.9 0
0
13
0 9 2 0 0 8192 0 0 11 9 0 3
428 304
428 315
486 315
13 1 3 0 0 4224 0 11 7 0 0 3
550 261
689 261
689 232
12 1 4 0 0 4224 0 11 8 0 0 3
550 270
731 270
731 253
11 1 5 0 0 4224 0 11 9 0 0 3
550 279
773 279
773 267
10 1 6 0 0 4224 0 11 10 0 0 3
550 288
811 288
811 283
0 8 7 0 0 12288 0 0 11 7 0 4
473 307
478 307
478 306
486 306
1 7 7 0 0 4224 0 1 11 0 0 4
374 331
473 331
473 297
486 297
0 6 2 0 0 0 0 0 11 9 0 3
478 288
478 288
486 288
1 5 2 0 0 4224 0 2 11 0 0 4
373 304
478 304
478 279
486 279
1 3 8 0 0 4224 0 4 11 0 0 4
375 257
478 257
478 261
486 261
1 4 9 0 0 4224 0 3 11 0 0 4
373 277
478 277
478 270
486 270
1 2 10 0 0 4224 0 5 11 0 0 4
374 229
473 229
473 252
486 252
1 1 11 0 0 4224 0 6 11 0 0 4
375 205
478 205
478 243
486 243
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
